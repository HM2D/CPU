`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:29:56 10/27/2015 
// Design Name: 
// Module Name:    MAINexp3 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module MAINexp3(clk,RD1,RD2,Output,Z
    );
	 input clk;
	 input [0:31] RD1,RD2;
	 output [0:31] Output;
	 output Z;
	 
	 MUX2_1 H1(R 
	 
	 
	 
	 


endmodule
